-- NO REGISTERS IN THIS STAGE, REGISTER FILE SAMPLES AT CLOCK EDGE ALREADY THUS IMPLEMENTING PIPELINE 
